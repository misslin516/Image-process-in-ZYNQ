`timescale 1ns / 1ps


module cos_table(
   input wire clk,
      
   input wire rd_en,
   input wire [8:0] addr,//0~360����ʾ��ת�Ƕ�
   
   output wire [8:0] dout
    );

    //��������
    reg [8:0] rom_data;
    
    //���
    always@(posedge clk ) begin
        if(rd_en) begin
            case(addr)
            default: rom_data <= 255;
            1: rom_data <= 254;
            2: rom_data <= 254;
            3: rom_data <= 254;
            4: rom_data <= 254;
            5: rom_data <= 254;
            6: rom_data <= 253;
            7: rom_data <= 253;
            8: rom_data <= 252;
            9: rom_data <= 251;
            10: rom_data <= 251;
            11: rom_data <= 250;
            12: rom_data <= 249;
            13: rom_data <= 248;
            14: rom_data <= 247;
            15: rom_data <= 246;
            16: rom_data <= 245;
            17: rom_data <= 243;
            18: rom_data <= 242;
            19: rom_data <= 241;
            20: rom_data <= 239;
            21: rom_data <= 238;
            22: rom_data <= 236;
            23: rom_data <= 234;
            24: rom_data <= 232;
            25: rom_data <= 231;
            26: rom_data <= 229;
            27: rom_data <= 227;
            28: rom_data <= 225;
            29: rom_data <= 223;
            30: rom_data <= 220;
            31: rom_data <= 218;
            32: rom_data <= 216;
            33: rom_data <= 213;
            34: rom_data <= 211;
            35: rom_data <= 208;
            36: rom_data <= 206;
            37: rom_data <= 203;
            38: rom_data <= 200;
            39: rom_data <= 198;
            40: rom_data <= 195;
            41: rom_data <= 192;
            42: rom_data <= 189;
            43: rom_data <= 186;
            44: rom_data <= 183;
            45: rom_data <= 180;
            46: rom_data <= 177;
            47: rom_data <= 173;
            48: rom_data <= 170;
            49: rom_data <= 167;
            50: rom_data <= 163;
            51: rom_data <= 160;
            52: rom_data <= 156;
            53: rom_data <= 153;
            54: rom_data <= 149;
            55: rom_data <= 146;
            56: rom_data <= 142;
            57: rom_data <= 138;
            58: rom_data <= 135;
            59: rom_data <= 131;
            60: rom_data <= 127;
            61: rom_data <= 123;
            62: rom_data <= 119;
            63: rom_data <= 115;
            64: rom_data <= 111;
            65: rom_data <= 107;
            66: rom_data <= 103;
            67: rom_data <= 99;
            68: rom_data <= 95;
            69: rom_data <= 91;
            70: rom_data <= 87;
            71: rom_data <= 83;
            72: rom_data <= 78;
            73: rom_data <= 74;
            74: rom_data <= 70;
            75: rom_data <= 65;
            76: rom_data <= 61;
            77: rom_data <= 57;
            78: rom_data <= 53;
            79: rom_data <= 48;
            80: rom_data <= 44;
            81: rom_data <= 39;
            82: rom_data <= 35;
            83: rom_data <= 31;
            84: rom_data <= 26;
            85: rom_data <= 22;
            86: rom_data <= 17;
            87: rom_data <= 13;
            88: rom_data <= 8;
            89: rom_data <= 4;
            90: rom_data <= 0;
            91: rom_data <= -4;
            92: rom_data <= -8;
            93: rom_data <= -13;
            94: rom_data <= -17;
            95: rom_data <= -22;
            96: rom_data <= -26;
            97: rom_data <= -31;
            98: rom_data <= -35;
            99: rom_data <= -39;
            100: rom_data <= -44;
            101: rom_data <= -48;
            102: rom_data <= -53;
            103: rom_data <= -57;
            104: rom_data <= -61;
            105: rom_data <= -65;
            106: rom_data <= -70;
            107: rom_data <= -74;
            108: rom_data <= -78;
            109: rom_data <= -83;
            110: rom_data <= -87;
            111: rom_data <= -91;
            112: rom_data <= -95;
            113: rom_data <= -99;
            114: rom_data <= -103;
            115: rom_data <= -107;
            116: rom_data <= -111;
            117: rom_data <= -115;
            118: rom_data <= -119;
            119: rom_data <= -123;
            120: rom_data <= -127;
            121: rom_data <= -131;
            122: rom_data <= -135;
            123: rom_data <= -138;
            124: rom_data <= -142;
            125: rom_data <= -146;
            126: rom_data <= -149;
            127: rom_data <= -153;
            128: rom_data <= -156;
            129: rom_data <= -160;
            130: rom_data <= -163;
            131: rom_data <= -167;
            132: rom_data <= -170;
            133: rom_data <= -173;
            134: rom_data <= -177;
            135: rom_data <= -180;
            136: rom_data <= -183;
            137: rom_data <= -186;
            138: rom_data <= -189;
            139: rom_data <= -192;
            140: rom_data <= -195;
            141: rom_data <= -198;
            142: rom_data <= -200;
            143: rom_data <= -203;
            144: rom_data <= -206;
            145: rom_data <= -208;
            146: rom_data <= -211;
            147: rom_data <= -213;
            148: rom_data <= -216;
            149: rom_data <= -218;
            150: rom_data <= -220;
            151: rom_data <= -223;
            152: rom_data <= -225;
            153: rom_data <= -227;
            154: rom_data <= -229;
            155: rom_data <= -231;
            156: rom_data <= -232;
            157: rom_data <= -234;
            158: rom_data <= -236;
            159: rom_data <= -238;
            160: rom_data <= -239;
            161: rom_data <= -241;
            162: rom_data <= -242;
            163: rom_data <= -243;
            164: rom_data <= -245;
            165: rom_data <= -246;
            166: rom_data <= -247;
            167: rom_data <= -248;
            168: rom_data <= -249;
            169: rom_data <= -250;
            170: rom_data <= -251;
            171: rom_data <= -251;
            172: rom_data <= -252;
            173: rom_data <= -253;
            174: rom_data <= -253;
            175: rom_data <= -254;
            176: rom_data <= -254;
            177: rom_data <= -254;
            178: rom_data <= -254;
            179: rom_data <= -254;
            180: rom_data <= -255;
            181: rom_data <= -254;
            182: rom_data <= -254;
            183: rom_data <= -254;
            184: rom_data <= -254;
            185: rom_data <= -254;
            186: rom_data <= -253;
            187: rom_data <= -253;
            188: rom_data <= -252;
            189: rom_data <= -251;
            190: rom_data <= -251;
            191: rom_data <= -250;
            192: rom_data <= -249;
            193: rom_data <= -248;
            194: rom_data <= -247;
            195: rom_data <= -246;
            196: rom_data <= -245;
            197: rom_data <= -243;
            198: rom_data <= -242;
            199: rom_data <= -241;
            200: rom_data <= -239;
            201: rom_data <= -238;
            202: rom_data <= -236;
            203: rom_data <= -234;
            204: rom_data <= -232;
            205: rom_data <= -231;
            206: rom_data <= -229;
            207: rom_data <= -227;
            208: rom_data <= -225;
            209: rom_data <= -223;
            210: rom_data <= -220;
            211: rom_data <= -218;
            212: rom_data <= -216;
            213: rom_data <= -213;
            214: rom_data <= -211;
            215: rom_data <= -208;
            216: rom_data <= -206;
            217: rom_data <= -203;
            218: rom_data <= -200;
            219: rom_data <= -198;
            220: rom_data <= -195;
            221: rom_data <= -192;
            222: rom_data <= -189;
            223: rom_data <= -186;
            224: rom_data <= -183;
            225: rom_data <= -180;
            226: rom_data <= -177;
            227: rom_data <= -173;
            228: rom_data <= -170;
            229: rom_data <= -167;
            230: rom_data <= -163;
            231: rom_data <= -160;
            232: rom_data <= -156;
            233: rom_data <= -153;
            234: rom_data <= -149;
            235: rom_data <= -146;
            236: rom_data <= -142;
            237: rom_data <= -138;
            238: rom_data <= -135;
            239: rom_data <= -131;
            240: rom_data <= -127;
            241: rom_data <= -123;
            242: rom_data <= -119;
            243: rom_data <= -115;
            244: rom_data <= -111;
            245: rom_data <= -107;
            246: rom_data <= -103;
            247: rom_data <= -99;
            248: rom_data <= -95;
            249: rom_data <= -91;
            250: rom_data <= -87;
            251: rom_data <= -83;
            252: rom_data <= -78;
            253: rom_data <= -74;
            254: rom_data <= -70;
            255: rom_data <= -65;
            256: rom_data <= -61;
            257: rom_data <= -57;
            258: rom_data <= -53;
            259: rom_data <= -48;
            260: rom_data <= -44;
            261: rom_data <= -39;
            262: rom_data <= -35;
            263: rom_data <= -31;
            264: rom_data <= -26;
            265: rom_data <= -22;
            266: rom_data <= -17;
            267: rom_data <= -13;
            268: rom_data <= -8;
            269: rom_data <= -4;
            270: rom_data <= 0;
            271: rom_data <= 4;
            272: rom_data <= 8;
            273: rom_data <= 13;
            274: rom_data <= 17;
            275: rom_data <= 22;
            276: rom_data <= 26;
            277: rom_data <= 31;
            278: rom_data <= 35;
            279: rom_data <= 39;
            280: rom_data <= 44;
            281: rom_data <= 48;
            282: rom_data <= 53;
            283: rom_data <= 57;
            284: rom_data <= 61;
            285: rom_data <= 65;
            286: rom_data <= 70;
            287: rom_data <= 74;
            288: rom_data <= 78;
            289: rom_data <= 83;
            290: rom_data <= 87;
            291: rom_data <= 91;
            292: rom_data <= 95;
            293: rom_data <= 99;
            294: rom_data <= 103;
            295: rom_data <= 107;
            296: rom_data <= 111;
            297: rom_data <= 115;
            298: rom_data <= 119;
            299: rom_data <= 123;
            300: rom_data <= 127;
            301: rom_data <= 131;
            302: rom_data <= 135;
            303: rom_data <= 138;
            304: rom_data <= 142;
            305: rom_data <= 146;
            306: rom_data <= 149;
            307: rom_data <= 153;
            308: rom_data <= 156;
            309: rom_data <= 160;
            310: rom_data <= 163;
            311: rom_data <= 167;
            312: rom_data <= 170;
            313: rom_data <= 173;
            314: rom_data <= 177;
            315: rom_data <= 180;
            316: rom_data <= 183;
            317: rom_data <= 186;
            318: rom_data <= 189;
            319: rom_data <= 192;
            320: rom_data <= 195;
            321: rom_data <= 198;
            322: rom_data <= 200;
            323: rom_data <= 203;
            324: rom_data <= 206;
            325: rom_data <= 208;
            326: rom_data <= 211;
            327: rom_data <= 213;
            328: rom_data <= 216;
            329: rom_data <= 218;
            330: rom_data <= 220;
            331: rom_data <= 223;
            332: rom_data <= 225;
            333: rom_data <= 227;
            334: rom_data <= 229;
            335: rom_data <= 231;
            336: rom_data <= 232;
            337: rom_data <= 234;
            338: rom_data <= 236;
            339: rom_data <= 238;
            340: rom_data <= 239;
            341: rom_data <= 241;
            342: rom_data <= 242;
            343: rom_data <= 243;
            344: rom_data <= 245;
            345: rom_data <= 246;
            346: rom_data <= 247;
            347: rom_data <= 248;
            348: rom_data <= 249;
            349: rom_data <= 250;
            350: rom_data <= 251;
            351: rom_data <= 251;
            352: rom_data <= 252;
            353: rom_data <= 253;
            354: rom_data <= 253;
            355: rom_data <= 254;
            356: rom_data <= 254;
            357: rom_data <= 254;
            358: rom_data <= 254;
            359: rom_data <= 254;            
            endcase
        end
    end
    
    assign dout = rom_data;
    
endmodule
